-- Copyright (C) 1991-2012 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 12.1 Build 243 01/31/2013 Service Pack 1 SJ Full Version"
-- CREATED		"Sun Aug 18 12:52:06 2013"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY controlBlock IS 
	PORT
	(
		SENSE_IN_HR :  IN  STD_LOGIC;
		SENSE_IN_VR :  IN  STD_LOGIC;
		CLK_IN :  IN  STD_LOGIC;
		PWM_IN_RIGHT :  IN  STD_LOGIC;
		SENSE_IN_HL :  IN  STD_LOGIC;
		PWM_IN_LEFT :  IN  STD_LOGIC;
		SENSE_IN_VL :  IN  STD_LOGIC;
		ABS_EN_GLOBAL :  IN  STD_LOGIC;
		PWM_OUT_VR :  OUT  STD_LOGIC;
		PWM_OUT_HR :  OUT  STD_LOGIC;
		OVERFLOW_LOW_OUT_HR :  OUT  STD_LOGIC;
		OVERFLOW_HIGH_OUT_HR :  OUT  STD_LOGIC;
		ABS_ENABLE_HR :  OUT  STD_LOGIC;
		BLOCK_DETECT_OUT_HR :  OUT  STD_LOGIC;
		PWM_OUT_HL :  OUT  STD_LOGIC;
		OVERFLOW_LOW_OUT_HL :  OUT  STD_LOGIC;
		OVERFLOW_HIGH_OUT_HL :  OUT  STD_LOGIC;
		ABS_ENABLE_HL :  OUT  STD_LOGIC;
		BLOCK_DETECT_OUT_HL :  OUT  STD_LOGIC;
		PWM_OUT_VL :  OUT  STD_LOGIC;
		OVERFLOW_LOW_OUT_VL :  OUT  STD_LOGIC;
		OVERFLOW_HIGH_OUT_VL :  OUT  STD_LOGIC;
		ABS_ENABLE_VL :  OUT  STD_LOGIC;
		BLOCK_DETECT_OUT_VL :  OUT  STD_LOGIC;
		OVERFLOW_LOW_OUT_VR :  OUT  STD_LOGIC;
		OVERFLOW_HIGH_OUT_VR :  OUT  STD_LOGIC;
		ABS_ENABLE_VR :  OUT  STD_LOGIC;
		BLOCK_DETECT_OUT_VR :  OUT  STD_LOGIC;
		LUT_INPUT_OUT :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		LUT_OUT :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		OUT_HIGH_HL :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		OUT_HIGH_HR :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		OUT_HIGH_VL :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		OUT_HIGH_VR :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		OUT_LOW_HL :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		OUT_LOW_HR :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		OUT_LOW_VL :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		OUT_LOW_VR :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END controlBlock;

ARCHITECTURE bdf_type OF controlBlock IS 

COMPONENT abscontrolhl
	PORT(CLK_IN : IN STD_LOGIC;
		 SENSE_IN_HL : IN STD_LOGIC;
		 PWM_IN_LEFT : IN STD_LOGIC;
		 ABS_EN_GLOBAL : IN STD_LOGIC;
		 COMPARATOR_SELECT_PORT_IN_HL : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 LUT_IN_HL : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 PWM_OUT_HL : OUT STD_LOGIC;
		 OVERFLOW_LOW_OUT_HL : OUT STD_LOGIC;
		 OVERFLOW_HIGH_OUT_HL : OUT STD_LOGIC;
		 ABS_ENABLE_OUT_HL : OUT STD_LOGIC;
		 BLOCK_DETECT_OUT_HL : OUT STD_LOGIC;
		 HIGH_LOW_MUX_OUT_HL : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 OUT_HIGH_HL : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 OUT_LOW_HL : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT abscontrolhr
	PORT(CLK_IN : IN STD_LOGIC;
		 SENSE_IN_HR : IN STD_LOGIC;
		 PWM_IN_RIGHT : IN STD_LOGIC;
		 ABS_EN_GLOBAL : IN STD_LOGIC;
		 COMPARATOR_SELECT_PORT_IN_HR : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 LUT_IN_HR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 PWM_OUT_HR : OUT STD_LOGIC;
		 OVERFLOW_LOW_OUT_HR : OUT STD_LOGIC;
		 OVERFLOW_HIGH_OUT_HR : OUT STD_LOGIC;
		 ABS_ENABLE_OUT_HR : OUT STD_LOGIC;
		 BLOCK_DETECT_OUT_HR : OUT STD_LOGIC;
		 HIGH_LOW_MUX_OUT_HR : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 OUT_HIGH_HR : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 OUT_LOW_HR : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT abscontrolvl
	PORT(CLK_IN : IN STD_LOGIC;
		 SENSE_IN_VL : IN STD_LOGIC;
		 PWM_IN_LEFT : IN STD_LOGIC;
		 ABS_EN_GLOBAL : IN STD_LOGIC;
		 COMPARATOR_SELECT_PORT_IN_VL : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 LUT_IN_VL : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 PWM_OUT_VL : OUT STD_LOGIC;
		 OVERFLOW_LOW_OUT_VL : OUT STD_LOGIC;
		 OVERFLOW_HIGH_OUT_VL : OUT STD_LOGIC;
		 ABS_ENABLE_OUT_VL : OUT STD_LOGIC;
		 BLOCK_DETECT_OUT_VL : OUT STD_LOGIC;
		 HIGH_LOW_MUX_OUT_VL : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 OUT_HIGH_VL : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 OUT_LOW_VL : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT abscontrolvr
	PORT(CLK_IN : IN STD_LOGIC;
		 SENSE_IN_VR : IN STD_LOGIC;
		 PWM_IN_RIGHT : IN STD_LOGIC;
		 ABS_EN_GLOBAL : IN STD_LOGIC;
		 COMPARATOR_SELECT_PORT_IN_VR : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 LUT_IN_VR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 PWM_OUT_VR : OUT STD_LOGIC;
		 OVERFLOW_LOW_OUT_VR : OUT STD_LOGIC;
		 OVERFLOW_HIGH_OUT_VR : OUT STD_LOGIC;
		 ABS_ENABLE_OUT_VR : OUT STD_LOGIC;
		 BLOCK_DETECT_OUT_VR : OUT STD_LOGIC;
		 HIGH_LOW_MUX_OUT_VR : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 OUT_HIGH_VR : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 OUT_LOW_VR : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lut
GENERIC (ADDR_WIDTH : INTEGER;
			DATA_WIDTH : INTEGER
			);
	PORT(clk : IN STD_LOGIC;
		 oldN : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 selectportin : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 maxN : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 selectportout : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lutmultiplexer
	PORT(clk : IN STD_LOGIC;
		 inport0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 inport1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 inport2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 inport3 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 outport : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 selectport : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	high_low_mux_out_hl :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	high_low_mux_out_hr :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	high_low_mux_out_vl :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	high_low_mux_out_vr :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	lut_out_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	lutmultiplexer_out :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	select_port :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC_VECTOR(1 DOWNTO 0);


BEGIN 



b2v_absControlHL_instance : abscontrolhl
PORT MAP(CLK_IN => CLK_IN,
		 SENSE_IN_HL => SENSE_IN_HL,
		 PWM_IN_LEFT => PWM_IN_LEFT,
		 ABS_EN_GLOBAL => ABS_EN_GLOBAL,
		 COMPARATOR_SELECT_PORT_IN_HL => select_port,
		 LUT_IN_HL => lut_out_ALTERA_SYNTHESIZED,
		 PWM_OUT_HL => PWM_OUT_HL,
		 OVERFLOW_LOW_OUT_HL => OVERFLOW_LOW_OUT_HL,
		 OVERFLOW_HIGH_OUT_HL => OVERFLOW_HIGH_OUT_HL,
		 ABS_ENABLE_OUT_HL => ABS_ENABLE_HL,
		 BLOCK_DETECT_OUT_HL => BLOCK_DETECT_OUT_HL,
		 HIGH_LOW_MUX_OUT_HL => high_low_mux_out_hl,
		 OUT_HIGH_HL => OUT_HIGH_HL,
		 OUT_LOW_HL => OUT_LOW_HL);


b2v_absControlHR_instance : abscontrolhr
PORT MAP(CLK_IN => CLK_IN,
		 SENSE_IN_HR => SENSE_IN_HR,
		 PWM_IN_RIGHT => PWM_IN_RIGHT,
		 ABS_EN_GLOBAL => ABS_EN_GLOBAL,
		 COMPARATOR_SELECT_PORT_IN_HR => select_port,
		 LUT_IN_HR => lut_out_ALTERA_SYNTHESIZED,
		 PWM_OUT_HR => PWM_OUT_HR,
		 OVERFLOW_LOW_OUT_HR => OVERFLOW_LOW_OUT_HR,
		 OVERFLOW_HIGH_OUT_HR => OVERFLOW_HIGH_OUT_HR,
		 ABS_ENABLE_OUT_HR => ABS_ENABLE_HR,
		 BLOCK_DETECT_OUT_HR => BLOCK_DETECT_OUT_HR,
		 HIGH_LOW_MUX_OUT_HR => high_low_mux_out_hr,
		 OUT_HIGH_HR => OUT_HIGH_HR,
		 OUT_LOW_HR => OUT_LOW_HR);


b2v_absControlVL_instance : abscontrolvl
PORT MAP(CLK_IN => CLK_IN,
		 SENSE_IN_VL => SENSE_IN_VL,
		 PWM_IN_LEFT => PWM_IN_LEFT,
		 ABS_EN_GLOBAL => ABS_EN_GLOBAL,
		 COMPARATOR_SELECT_PORT_IN_VL => select_port,
		 LUT_IN_VL => lut_out_ALTERA_SYNTHESIZED,
		 PWM_OUT_VL => PWM_OUT_VL,
		 OVERFLOW_LOW_OUT_VL => OVERFLOW_LOW_OUT_VL,
		 OVERFLOW_HIGH_OUT_VL => OVERFLOW_HIGH_OUT_VL,
		 ABS_ENABLE_OUT_VL => ABS_ENABLE_VL,
		 BLOCK_DETECT_OUT_VL => BLOCK_DETECT_OUT_VL,
		 HIGH_LOW_MUX_OUT_VL => high_low_mux_out_vl,
		 OUT_HIGH_VL => OUT_HIGH_VL,
		 OUT_LOW_VL => OUT_LOW_VL);


b2v_absControlVR_instance : abscontrolvr
PORT MAP(CLK_IN => CLK_IN,
		 SENSE_IN_VR => SENSE_IN_VR,
		 PWM_IN_RIGHT => PWM_IN_RIGHT,
		 ABS_EN_GLOBAL => ABS_EN_GLOBAL,
		 COMPARATOR_SELECT_PORT_IN_VR => select_port,
		 LUT_IN_VR => lut_out_ALTERA_SYNTHESIZED,
		 PWM_OUT_VR => PWM_OUT_VR,
		 OVERFLOW_LOW_OUT_VR => OVERFLOW_LOW_OUT_VR,
		 OVERFLOW_HIGH_OUT_VR => OVERFLOW_HIGH_OUT_VR,
		 ABS_ENABLE_OUT_VR => ABS_ENABLE_VR,
		 BLOCK_DETECT_OUT_VR => BLOCK_DETECT_OUT_VR,
		 HIGH_LOW_MUX_OUT_VR => high_low_mux_out_vr,
		 OUT_HIGH_VR => OUT_HIGH_VR,
		 OUT_LOW_VR => OUT_LOW_VR);


b2v_inst3 : lut
GENERIC MAP(ADDR_WIDTH => 14,
			DATA_WIDTH => 16
			)
PORT MAP(clk => CLK_IN,
		 oldN => lutmultiplexer_out(13 DOWNTO 0),
		 selectportin => SYNTHESIZED_WIRE_0,
		 maxN => lut_out_ALTERA_SYNTHESIZED,
		 selectportout => select_port);


b2v_lutmultiplexer : lutmultiplexer
PORT MAP(clk => CLK_IN,
		 inport0 => high_low_mux_out_hr,
		 inport1 => high_low_mux_out_vr,
		 inport2 => high_low_mux_out_hl,
		 inport3 => high_low_mux_out_vl,
		 outport => lutmultiplexer_out,
		 selectport => SYNTHESIZED_WIRE_0);

LUT_INPUT_OUT <= lutmultiplexer_out;
LUT_OUT <= lut_out_ALTERA_SYNTHESIZED;

END bdf_type;